../../Tiny_TCM/fabrics/AHBL/src_tb/AHBL_Target_AXI4_Initiator.bsv